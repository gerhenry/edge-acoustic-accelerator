* Placeholder ngspice testbench
.end
