// Stub RTL
module user_regbank(); endmodule
