* Include your PDK models here
